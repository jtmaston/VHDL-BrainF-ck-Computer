library ieee;
use ieee.std_logic_1164.all;

package bfCPUDataTypes is
    type addressBus is array(0 to 7) of std_logic;
end bfCPUDataTypes;